    // // Parameters for burst types
    // parameter single = 3'b000;
    // parameter incr   = 3'b001;
    // parameter wrap4  = 3'b010;
    // parameter incr4  = 3'b011;
    // parameter wrap8  = 3'b100;
    // parameter incr8  = 3'b101;
    // parameter wrap16 = 3'b110;
    // parameter incr16 = 3'b111;

    //     // Task to get address
    //     task get_address(output bit [31:0] addr);
    //         wait(ahb_vif.HREADY);
    //         addr = ahb_vif.HADDR;
    //     endtask